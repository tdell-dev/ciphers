module simon_enc_subkey #( ) (
	input clk,
	input rst,
	input [255:0] enc_key_in,
	input         enc_key_in_vld,
	output        enc_key_in_rdy
);

    wire clk;
    wire rst;
    wire [255:0] enc_key_in;
    wire enc_key_in_vld;
    reg  enc_key_in_rdy;



endmodule

